module HazardUnit
(
input [4:0] Instruction_ID,
input [4:0] MemRead_EX,
input [4:0] RT_EX,
output [1:0] DWrite,
output [1:0] PCWrite,
output [1:0] Hazardflush

);

endmodule
