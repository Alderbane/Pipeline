/******************************************************************
* Description
*		This is the HazardUnit:
* Version:
*	1.0
* Author:
*Luis David Gallegos Godoy
* email:
*	is709571@iteso.mx
* Date:
*	17/07/2019
******************************************************************/
module Hazard
(
input [4:0] Instruction_ID,
input [4:0] RT_EX,
input MemRead_EX,
output DWrite,
output PCWrite,
output Bubble

);

endmodule
